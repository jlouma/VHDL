----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:47:08 01/25/2015 
-- Design Name: 
-- Module Name:    BaudCLKGen - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BaudCLKGen is
    Port ( BaudSel : in  STD_LOGIC_VECTOR (2 downto 0);
           CLK : in  STD_LOGIC;
           BaudCLK : out  STD_LOGIC);
end BaudCLKGen;

architecture Behavioral of BaudCLKGen is

begin


end Behavioral;

